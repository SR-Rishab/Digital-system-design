module mux16_tb();
wire y;
reg  [3:0]s;
reg [15:0]d;
mux16 m0(s,d,y);
initial
begin
d = 16'b1010_1010_1010_1010;
s = 4'b0000;
#10;
d = 16'b1010_1010_1010_1010;
s = 4'b0001;
#10;
d = 16'b1010_1010_1010_1010;
s = 4'b0010;
#10;
d = 16'b1010_1010_1010_1010;
s = 4'b0011;
#10;
end
endmodule
